`timescale 1ns / 1ps
//~ ////////////////////////////////////////////////////////////////////////////////
//! Company: Bug Makers Inc.
//! Engineer:  👽
//~ 
//! Create Date:    19:12:12 10/16/2025
//! Design Name:
//! Module Name:    main_memory
//! Project Name: 🐞

//~ ///////////////////////////////////////////////////////////////////////////////////////////////



module main_memory(
    input wire clk,
    input wire reset,
    
)